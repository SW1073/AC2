--
-- Copyright (c) 2018, UPC
-- All rights reserved.
-- 

library ieee;
use ieee.std_logic_1164.all;

use work.cte_tipos_deco_camino_pkg.all;
use work.componentes_control_seg_pkg.all;
use work.retardos_cntl_seg_pkg.all;

entity LDRS is
	port(opsecDL, opsecA : in st_opSEC;
		RS: out std_logic);
end LDRS;


architecture comportamiento of LDRS is

begin

	RS <= (opsecDL(num_opSEC-1) or opsecA(num_opSEC-1)) after retLDRS;
	
end comportamiento;
